--UserModule_Simulation_Waveform1.vhdl
--
--SpaceWire Board / User FPGA / Modularized Structure Template
--UserFPGA Simulation / sample waveform generator
--
--ver20071128 Takayuki Yuasa
--file created

---------------------------------------------------
--Declarations of Libraries
---------------------------------------------------
library ieee,work;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.iBus_Library.all;
use work.iBus_AddressMap.all;
use work.UserModule_Library.all;

---------------------------------------------------
--Entity Declaration
---------------------------------------------------
entity UserModule_Simulation_Waveform1 is
	port(
		Start		:	in	std_logic;
		waveform	:	out std_logic_vector(15 downto 0);
		--clock and reset
		Clock			:	in		std_logic;
		GlobalReset	:	in		std_logic
	);
end UserModule_Simulation_Waveform1;

---------------------------------------------------
--Behavioral description
---------------------------------------------------
architecture Behavioral of UserModule_Simulation_Waveform1 is

	---------------------------------------------------
	--Declarations of Components
	---------------------------------------------------

	---------------------------------------------------
	--Declarations of Signals
	---------------------------------------------------
	
	signal flag : std_logic := '0';
	type vector16 is array (INTEGER range <>) of std_logic_vector(15 downto 0);
	signal wave : vector16(800 downto 0);
	signal i : integer :=0;
	--Registers

	---------------------------------------------------
	--Beginning of behavioral description
	---------------------------------------------------
	begin	
	
	---------------------------------------------------
	--Instantiations of Components
	---------------------------------------------------

	---------------------------------------------------
	--Static relationships
	---------------------------------------------------
	waveform <= wave(i);
	
	---------------------------------------------------
	--Dynamic Processes with Sensitivity List
	---------------------------------------------------

	process (Clock, GlobalReset)
	begin
		if (GlobalReset='0') then
			i <= 0;
		elsif (Clock'Event and Clock='1') then
			if (flag='1') then
				if (i<750) then
					i <= i + 1;
				end if;
			else
				if (start='1') then
					flag <= '1';
				end if;
			end if;
		end if;
	end process;
	
	wave(0) <= conv_std_logic_vector(1,16);
	wave(1) <= conv_std_logic_vector(2,16);
	wave(2) <= conv_std_logic_vector(3,16);
	wave(3) <= conv_std_logic_vector(4,16);
	wave(4) <= conv_std_logic_vector(5,16);
	wave(5) <= conv_std_logic_vector(6,16);
	wave(6) <= conv_std_logic_vector(7,16);
	wave(7) <= conv_std_logic_vector(8,16);
	wave(8) <= conv_std_logic_vector(9,16);
	wave(9) <= conv_std_logic_vector(2039,16);
	wave(10) <= conv_std_logic_vector(2028,16);
	wave(11) <= conv_std_logic_vector(2052,16);
	wave(12) <= conv_std_logic_vector(2069,16);
	wave(13) <= conv_std_logic_vector(2063,16);
	wave(14) <= conv_std_logic_vector(2064,16);
	wave(15) <= conv_std_logic_vector(2106,16);
	wave(16) <= conv_std_logic_vector(2170,16);
	wave(17) <= conv_std_logic_vector(2224,16);
	wave(18) <= conv_std_logic_vector(2285,16);
	wave(19) <= conv_std_logic_vector(2377,16);
	wave(20) <= conv_std_logic_vector(2490,16);
	wave(21) <= conv_std_logic_vector(2603,16);
	wave(22) <= conv_std_logic_vector(2717,16);
	wave(23) <= conv_std_logic_vector(2840,16);
	wave(24) <= conv_std_logic_vector(2963,16);
	wave(25) <= conv_std_logic_vector(3082,16);
	wave(26) <= conv_std_logic_vector(3194,16);
	wave(27) <= conv_std_logic_vector(3296,16);
	wave(28) <= conv_std_logic_vector(3385,16);
	wave(29) <= conv_std_logic_vector(3462,16);
	wave(30) <= conv_std_logic_vector(3521,16);
	wave(31) <= conv_std_logic_vector(3564,16);
	wave(32) <= conv_std_logic_vector(3590,16);
	wave(33) <= conv_std_logic_vector(3599,16);
	wave(34) <= conv_std_logic_vector(3592,16);
	wave(35) <= conv_std_logic_vector(3568,16);
	wave(36) <= conv_std_logic_vector(3531,16);
	wave(37) <= conv_std_logic_vector(3480,16);
	wave(38) <= conv_std_logic_vector(3417,16);
	wave(39) <= conv_std_logic_vector(3345,16);
	wave(40) <= conv_std_logic_vector(3264,16);
	wave(41) <= conv_std_logic_vector(3177,16);
	wave(42) <= conv_std_logic_vector(3085,16);
	wave(43) <= conv_std_logic_vector(2990,16);
	wave(44) <= conv_std_logic_vector(2894,16);
	wave(45) <= conv_std_logic_vector(2797,16);
	wave(46) <= conv_std_logic_vector(2702,16);
	wave(47) <= conv_std_logic_vector(2607,16);
	wave(48) <= conv_std_logic_vector(2517,16);
	wave(49) <= conv_std_logic_vector(2430,16);
	wave(50) <= conv_std_logic_vector(2347,16);
	wave(51) <= conv_std_logic_vector(2269,16);
	wave(52) <= conv_std_logic_vector(2197,16);
	wave(53) <= conv_std_logic_vector(2131,16);
	wave(54) <= conv_std_logic_vector(2065,16);
	wave(55) <= conv_std_logic_vector(2005,16);
	wave(56) <= conv_std_logic_vector(1959,16);
	wave(57) <= conv_std_logic_vector(1921,16);
	wave(58) <= conv_std_logic_vector(1877,16);
	wave(59) <= conv_std_logic_vector(1824,16);
	wave(60) <= conv_std_logic_vector(1789,16);
	wave(61) <= conv_std_logic_vector(1789,16);
	wave(62) <= conv_std_logic_vector(1774,16);
	wave(63) <= conv_std_logic_vector(1718,16);
	wave(64) <= conv_std_logic_vector(1688,16);
	wave(65) <= conv_std_logic_vector(1709,16);
	wave(66) <= conv_std_logic_vector(1711,16);
	wave(67) <= conv_std_logic_vector(1663,16);
	wave(68) <= conv_std_logic_vector(1639,16);
	wave(69) <= conv_std_logic_vector(1669,16);
	wave(70) <= conv_std_logic_vector(1683,16);
	wave(71) <= conv_std_logic_vector(1644,16);
	wave(72) <= conv_std_logic_vector(1620,16);
	wave(73) <= conv_std_logic_vector(1653,16);
	wave(74) <= conv_std_logic_vector(1674,16);
	wave(75) <= conv_std_logic_vector(1644,16);
	wave(76) <= conv_std_logic_vector(1619,16);
	wave(77) <= conv_std_logic_vector(1651,16);
	wave(78) <= conv_std_logic_vector(1679,16);
	wave(79) <= conv_std_logic_vector(1654,16);
	wave(80) <= conv_std_logic_vector(1627,16);
	wave(81) <= conv_std_logic_vector(1656,16);
	wave(82) <= conv_std_logic_vector(1691,16);
	wave(83) <= conv_std_logic_vector(1670,16);
	wave(84) <= conv_std_logic_vector(1640,16);
	wave(85) <= conv_std_logic_vector(1666,16);
	wave(86) <= conv_std_logic_vector(1702,16);
	wave(87) <= conv_std_logic_vector(1689,16);
	wave(88) <= conv_std_logic_vector(1658,16);
	wave(89) <= conv_std_logic_vector(1676,16);
	wave(90) <= conv_std_logic_vector(1716,16);
	wave(91) <= conv_std_logic_vector(1711,16);
	wave(92) <= conv_std_logic_vector(1679,16);
	wave(93) <= conv_std_logic_vector(1687,16);
	wave(94) <= conv_std_logic_vector(1728,16);
	wave(95) <= conv_std_logic_vector(1735,16);
	wave(96) <= conv_std_logic_vector(1701,16);
	wave(97) <= conv_std_logic_vector(1700,16);
	wave(98) <= conv_std_logic_vector(1741,16);
	wave(99) <= conv_std_logic_vector(1754,16);
	wave(100) <= conv_std_logic_vector(1722,16);
	wave(101) <= conv_std_logic_vector(1715,16);
	wave(102) <= conv_std_logic_vector(1752,16);
	wave(103) <= conv_std_logic_vector(1769,16);
	wave(104) <= conv_std_logic_vector(1746,16);
	wave(105) <= conv_std_logic_vector(1730,16);
	wave(106) <= conv_std_logic_vector(1761,16);
	wave(107) <= conv_std_logic_vector(1789,16);
	wave(108) <= conv_std_logic_vector(1769,16);
	wave(109) <= conv_std_logic_vector(1745,16);
	wave(110) <= conv_std_logic_vector(1770,16);
	wave(111) <= conv_std_logic_vector(1805,16);
	wave(112) <= conv_std_logic_vector(1790,16);
	wave(113) <= conv_std_logic_vector(1761,16);
	wave(114) <= conv_std_logic_vector(1780,16);
	wave(115) <= conv_std_logic_vector(1815,16);
	wave(116) <= conv_std_logic_vector(1810,16);
	wave(117) <= conv_std_logic_vector(1780,16);
	wave(118) <= conv_std_logic_vector(1788,16);
	wave(119) <= conv_std_logic_vector(1824,16);
	wave(120) <= conv_std_logic_vector(1829,16);
	wave(121) <= conv_std_logic_vector(1797,16);
	wave(122) <= conv_std_logic_vector(1798,16);
	wave(123) <= conv_std_logic_vector(1837,16);
	wave(124) <= conv_std_logic_vector(1847,16);
	wave(125) <= conv_std_logic_vector(1816,16);
	wave(126) <= conv_std_logic_vector(1807,16);
	wave(127) <= conv_std_logic_vector(1844,16);
	wave(128) <= conv_std_logic_vector(1860,16);
	wave(129) <= conv_std_logic_vector(1835,16);
	wave(130) <= conv_std_logic_vector(1819,16);
	wave(131) <= conv_std_logic_vector(1848,16);
	wave(132) <= conv_std_logic_vector(1873,16);
	wave(133) <= conv_std_logic_vector(1852,16);
	wave(134) <= conv_std_logic_vector(1831,16);
	wave(135) <= conv_std_logic_vector(1855,16);
	wave(136) <= conv_std_logic_vector(1883,16);
	wave(137) <= conv_std_logic_vector(1871,16);
	wave(138) <= conv_std_logic_vector(1844,16);
	wave(139) <= conv_std_logic_vector(1859,16);
	wave(140) <= conv_std_logic_vector(1893,16);
	wave(141) <= conv_std_logic_vector(1888,16);
	wave(142) <= conv_std_logic_vector(1859,16);
	wave(143) <= conv_std_logic_vector(1864,16);
	wave(144) <= conv_std_logic_vector(1900,16);
	wave(145) <= conv_std_logic_vector(1905,16);
	wave(146) <= conv_std_logic_vector(1873,16);
	wave(147) <= conv_std_logic_vector(1870,16);
	wave(148) <= conv_std_logic_vector(1906,16);
	wave(149) <= conv_std_logic_vector(1917,16);
	wave(150) <= conv_std_logic_vector(1891,16);
	wave(151) <= conv_std_logic_vector(1876,16);
	wave(152) <= conv_std_logic_vector(1907,16);
	wave(153) <= conv_std_logic_vector(1929,16);
	wave(154) <= conv_std_logic_vector(1908,16);
	wave(155) <= conv_std_logic_vector(1887,16);
	wave(156) <= conv_std_logic_vector(1908,16);
	wave(157) <= conv_std_logic_vector(1936,16);
	wave(158) <= conv_std_logic_vector(1925,16);
	wave(159) <= conv_std_logic_vector(1897,16);
	wave(160) <= conv_std_logic_vector(1912,16);
	wave(161) <= conv_std_logic_vector(1943,16);
	wave(162) <= conv_std_logic_vector(1938,16);
	wave(163) <= conv_std_logic_vector(1910,16);
	wave(164) <= conv_std_logic_vector(1914,16);
	wave(165) <= conv_std_logic_vector(1946,16);
	wave(166) <= conv_std_logic_vector(1952,16);
	wave(167) <= conv_std_logic_vector(1923,16);
	wave(168) <= conv_std_logic_vector(1917,16);
	wave(169) <= conv_std_logic_vector(1949,16);
	wave(170) <= conv_std_logic_vector(1961,16);
	wave(171) <= conv_std_logic_vector(1936,16);
	wave(172) <= conv_std_logic_vector(1923,16);
	wave(173) <= conv_std_logic_vector(1948,16);
	wave(174) <= conv_std_logic_vector(1969,16);
	wave(175) <= conv_std_logic_vector(1951,16);
	wave(176) <= conv_std_logic_vector(1929,16);
	wave(177) <= conv_std_logic_vector(1947,16);
	wave(178) <= conv_std_logic_vector(1974,16);
	wave(179) <= conv_std_logic_vector(1964,16);
	wave(180) <= conv_std_logic_vector(1937,16);
	wave(181) <= conv_std_logic_vector(1948,16);
	wave(182) <= conv_std_logic_vector(1977,16);
	wave(183) <= conv_std_logic_vector(1976,16);
	wave(184) <= conv_std_logic_vector(1949,16);
	wave(185) <= conv_std_logic_vector(1948,16);
	wave(186) <= conv_std_logic_vector(1977,16);
	wave(187) <= conv_std_logic_vector(1987,16);
	wave(188) <= conv_std_logic_vector(1960,16);
	wave(189) <= conv_std_logic_vector(1949,16);
	wave(190) <= conv_std_logic_vector(1977,16);
	wave(191) <= conv_std_logic_vector(1992,16);
	wave(192) <= conv_std_logic_vector(1974,16);
	wave(193) <= conv_std_logic_vector(1955,16);
	wave(194) <= conv_std_logic_vector(1971,16);
	wave(195) <= conv_std_logic_vector(1996,16);
	wave(196) <= conv_std_logic_vector(1989,16);
	wave(197) <= conv_std_logic_vector(1964,16);
	wave(198) <= conv_std_logic_vector(1968,16);
	wave(199) <= conv_std_logic_vector(1998,16);
	wave(200) <= conv_std_logic_vector(2001,16);
	wave(201) <= conv_std_logic_vector(1973,16);
	wave(202) <= conv_std_logic_vector(1968,16);
	wave(203) <= conv_std_logic_vector(1998,16);
	wave(204) <= conv_std_logic_vector(2008,16);
	wave(205) <= conv_std_logic_vector(1981,16);
	wave(206) <= conv_std_logic_vector(1971,16);
	wave(207) <= conv_std_logic_vector(1998,16);
	wave(208) <= conv_std_logic_vector(2015,16);
	wave(209) <= conv_std_logic_vector(1995,16);
	wave(210) <= conv_std_logic_vector(1975,16);
	wave(211) <= conv_std_logic_vector(1993,16);
	wave(212) <= conv_std_logic_vector(2015,16);
	wave(213) <= conv_std_logic_vector(2003,16);
	wave(214) <= conv_std_logic_vector(1981,16);
	wave(215) <= conv_std_logic_vector(1991,16);
	wave(216) <= conv_std_logic_vector(2018,16);
	wave(217) <= conv_std_logic_vector(2015,16);
	wave(218) <= conv_std_logic_vector(1988,16);
	wave(219) <= conv_std_logic_vector(1989,16);
	wave(220) <= conv_std_logic_vector(2017,16);
	wave(221) <= conv_std_logic_vector(2023,16);
	wave(222) <= conv_std_logic_vector(1998,16);
	wave(223) <= conv_std_logic_vector(1988,16);
	wave(224) <= conv_std_logic_vector(2015,16);
	wave(225) <= conv_std_logic_vector(2029,16);
	wave(226) <= conv_std_logic_vector(2007,16);
	wave(227) <= conv_std_logic_vector(1990,16);
	wave(228) <= conv_std_logic_vector(2011,16);
	wave(229) <= conv_std_logic_vector(2033,16);
	wave(230) <= conv_std_logic_vector(2017,16);
	wave(231) <= conv_std_logic_vector(1994,16);
	wave(232) <= conv_std_logic_vector(2007,16);
	wave(233) <= conv_std_logic_vector(2033,16);
	wave(234) <= conv_std_logic_vector(2026,16);
	wave(235) <= conv_std_logic_vector(2000,16);
	wave(236) <= conv_std_logic_vector(2003,16);
	wave(237) <= conv_std_logic_vector(2032,16);
	wave(238) <= conv_std_logic_vector(2034,16);
	wave(239) <= conv_std_logic_vector(2008,16);
	wave(240) <= conv_std_logic_vector(2002,16);
	wave(241) <= conv_std_logic_vector(2029,16);
	wave(242) <= conv_std_logic_vector(2041,16);
	wave(243) <= conv_std_logic_vector(2017,16);
	wave(244) <= conv_std_logic_vector(2002,16);
	wave(245) <= conv_std_logic_vector(2024,16);
	wave(246) <= conv_std_logic_vector(2044,16);
	wave(247) <= conv_std_logic_vector(2026,16);
	wave(248) <= conv_std_logic_vector(2005,16);
	wave(249) <= conv_std_logic_vector(2019,16);
	wave(250) <= conv_std_logic_vector(2043,16);
	wave(251) <= conv_std_logic_vector(2036,16);
	wave(252) <= conv_std_logic_vector(2012,16);
	wave(253) <= conv_std_logic_vector(2014,16);
	wave(254) <= conv_std_logic_vector(2041,16);
	wave(255) <= conv_std_logic_vector(2045,16);
	wave(256) <= conv_std_logic_vector(2019,16);
	wave(257) <= conv_std_logic_vector(2012,16);
	wave(258) <= conv_std_logic_vector(2037,16);
	wave(259) <= conv_std_logic_vector(2049,16);
	wave(260) <= conv_std_logic_vector(2029,16);
	wave(261) <= conv_std_logic_vector(2012,16);
	wave(262) <= conv_std_logic_vector(2032,16);
	wave(263) <= conv_std_logic_vector(2052,16);
	wave(264) <= conv_std_logic_vector(2038,16);
	wave(265) <= conv_std_logic_vector(2014,16);
	wave(266) <= conv_std_logic_vector(2027,16);
	wave(267) <= conv_std_logic_vector(2053,16);
	wave(268) <= conv_std_logic_vector(2046,16);
	wave(269) <= conv_std_logic_vector(2019,16);
	wave(270) <= conv_std_logic_vector(2023,16);
	wave(271) <= conv_std_logic_vector(2050,16);
	wave(272) <= conv_std_logic_vector(2053,16);
	wave(273) <= conv_std_logic_vector(2027,16);
	wave(274) <= conv_std_logic_vector(2020,16);
	wave(275) <= conv_std_logic_vector(2045,16);
	wave(276) <= conv_std_logic_vector(2057,16);
	wave(277) <= conv_std_logic_vector(2035,16);
	wave(278) <= conv_std_logic_vector(2019,16);
	wave(279) <= conv_std_logic_vector(2040,16);
	wave(280) <= conv_std_logic_vector(2060,16);
	wave(281) <= conv_std_logic_vector(2043,16);
	wave(282) <= conv_std_logic_vector(2018,16);
	wave(283) <= conv_std_logic_vector(2038,16);
	wave(284) <= conv_std_logic_vector(2062,16);
	wave(285) <= conv_std_logic_vector(2045,16);
	wave(286) <= conv_std_logic_vector(2021,16);
	wave(287) <= conv_std_logic_vector(2035,16);
	wave(288) <= conv_std_logic_vector(2060,16);
	wave(289) <= conv_std_logic_vector(2053,16);
	wave(290) <= conv_std_logic_vector(2027,16);
	wave(291) <= conv_std_logic_vector(2030,16);
	wave(292) <= conv_std_logic_vector(2057,16);
	wave(293) <= conv_std_logic_vector(2059,16);
	wave(294) <= conv_std_logic_vector(2033,16);
	wave(295) <= conv_std_logic_vector(2026,16);
	wave(296) <= conv_std_logic_vector(2052,16);
	wave(297) <= conv_std_logic_vector(2062,16);
	wave(298) <= conv_std_logic_vector(2038,16);
	wave(299) <= conv_std_logic_vector(2025,16);
	wave(300) <= conv_std_logic_vector(2047,16);
	wave(301) <= conv_std_logic_vector(2066,16);
	wave(302) <= conv_std_logic_vector(2049,16);
	wave(303) <= conv_std_logic_vector(2028,16);
	wave(304) <= conv_std_logic_vector(2039,16);
	wave(305) <= conv_std_logic_vector(2062,16);
	wave(306) <= conv_std_logic_vector(2057,16);
	wave(307) <= conv_std_logic_vector(2031,16);
	wave(308) <= conv_std_logic_vector(2033,16);
	wave(309) <= conv_std_logic_vector(2059,16);
	wave(310) <= conv_std_logic_vector(2063,16);
	wave(311) <= conv_std_logic_vector(2038,16);
	wave(312) <= conv_std_logic_vector(2029,16);
	wave(313) <= conv_std_logic_vector(2054,16);
	wave(314) <= conv_std_logic_vector(2067,16);
	wave(315) <= conv_std_logic_vector(2045,16);
	wave(316) <= conv_std_logic_vector(2028,16);
	wave(317) <= conv_std_logic_vector(2049,16);
	wave(318) <= conv_std_logic_vector(2067,16);
	wave(319) <= conv_std_logic_vector(2050,16);
	wave(320) <= conv_std_logic_vector(2028,16);
	wave(321) <= conv_std_logic_vector(2044,16);
	wave(322) <= conv_std_logic_vector(2067,16);
	wave(323) <= conv_std_logic_vector(2056,16);
	wave(324) <= conv_std_logic_vector(2031,16);
	wave(325) <= conv_std_logic_vector(2038,16);
	wave(326) <= conv_std_logic_vector(2065,16);
	wave(327) <= conv_std_logic_vector(2062,16);
	wave(328) <= conv_std_logic_vector(2035,16);
	wave(329) <= conv_std_logic_vector(2034,16);
	wave(330) <= conv_std_logic_vector(2059,16);
	wave(331) <= conv_std_logic_vector(2066,16);
	wave(332) <= conv_std_logic_vector(2042,16);
	wave(333) <= conv_std_logic_vector(2030,16);
	wave(334) <= conv_std_logic_vector(2053,16);
	wave(335) <= conv_std_logic_vector(2068,16);
	wave(336) <= conv_std_logic_vector(2048,16);
	wave(337) <= conv_std_logic_vector(2029,16);
	wave(338) <= conv_std_logic_vector(2047,16);
	wave(339) <= conv_std_logic_vector(2068,16);
	wave(340) <= conv_std_logic_vector(2055,16);
	wave(341) <= conv_std_logic_vector(2032,16);
	wave(342) <= conv_std_logic_vector(2040,16);
	wave(343) <= conv_std_logic_vector(2065,16);
	wave(344) <= conv_std_logic_vector(2062,16);
	wave(345) <= conv_std_logic_vector(2036,16);
	wave(346) <= conv_std_logic_vector(2034,16);
	wave(347) <= conv_std_logic_vector(2062,16);
	wave(348) <= conv_std_logic_vector(2067,16);
	wave(349) <= conv_std_logic_vector(2041,16);
	wave(350) <= conv_std_logic_vector(2032,16);
	wave(351) <= conv_std_logic_vector(2057,16);
	wave(352) <= conv_std_logic_vector(2070,16);
	wave(353) <= conv_std_logic_vector(2048,16);
	wave(354) <= conv_std_logic_vector(2032,16);
	wave(355) <= conv_std_logic_vector(2052,16);
	wave(356) <= conv_std_logic_vector(2071,16);
	wave(357) <= conv_std_logic_vector(2055,16);
	wave(358) <= conv_std_logic_vector(2033,16);
	wave(359) <= conv_std_logic_vector(2046,16);
	wave(360) <= conv_std_logic_vector(2069,16);
	wave(361) <= conv_std_logic_vector(2063,16);
	wave(362) <= conv_std_logic_vector(2036,16);
	wave(363) <= conv_std_logic_vector(2040,16);
	wave(364) <= conv_std_logic_vector(2066,16);
	wave(365) <= conv_std_logic_vector(2068,16);
	wave(366) <= conv_std_logic_vector(2042,16);
	wave(367) <= conv_std_logic_vector(2035,16);
	wave(368) <= conv_std_logic_vector(2061,16);
	wave(369) <= conv_std_logic_vector(2071,16);
	wave(370) <= conv_std_logic_vector(2048,16);
	wave(371) <= conv_std_logic_vector(2036,16);
	wave(372) <= conv_std_logic_vector(2054,16);
	wave(373) <= conv_std_logic_vector(2068,16);
	wave(374) <= conv_std_logic_vector(2057,16);
	wave(375) <= conv_std_logic_vector(2036,16);
	wave(376) <= conv_std_logic_vector(2043,16);
	wave(377) <= conv_std_logic_vector(2067,16);
	wave(378) <= conv_std_logic_vector(2066,16);
	wave(379) <= conv_std_logic_vector(2039,16);
	wave(380) <= conv_std_logic_vector(2037,16);
	wave(381) <= conv_std_logic_vector(2063,16);
	wave(382) <= conv_std_logic_vector(2070,16);
	wave(383) <= conv_std_logic_vector(2044,16);
	wave(384) <= conv_std_logic_vector(2034,16);
	wave(385) <= conv_std_logic_vector(2058,16);
	wave(386) <= conv_std_logic_vector(2071,16);
	wave(387) <= conv_std_logic_vector(2051,16);
	wave(388) <= conv_std_logic_vector(2036,16);
	wave(389) <= conv_std_logic_vector(2050,16);
	wave(390) <= conv_std_logic_vector(2072,16);
	wave(391) <= conv_std_logic_vector(2059,16);
	wave(392) <= conv_std_logic_vector(2033,16);
	wave(393) <= conv_std_logic_vector(2045,16);
	wave(394) <= conv_std_logic_vector(2069,16);
	wave(395) <= conv_std_logic_vector(2064,16);
	wave(396) <= conv_std_logic_vector(2040,16);
	wave(397) <= conv_std_logic_vector(2035,16);
	wave(398) <= conv_std_logic_vector(2066,16);
	wave(399) <= conv_std_logic_vector(2068,16);
	wave(400) <= conv_std_logic_vector(2045,16);
	wave(401) <= conv_std_logic_vector(2036,16);
	wave(402) <= conv_std_logic_vector(2053,16);
	wave(403) <= conv_std_logic_vector(2072,16);
	wave(404) <= conv_std_logic_vector(2055,16);
	wave(405) <= conv_std_logic_vector(2032,16);
	wave(406) <= conv_std_logic_vector(2047,16);
	wave(407) <= conv_std_logic_vector(2071,16);
	wave(408) <= conv_std_logic_vector(2060,16);
	wave(409) <= conv_std_logic_vector(2036,16);
	wave(410) <= conv_std_logic_vector(2041,16);
	wave(411) <= conv_std_logic_vector(2066,16);
	wave(412) <= conv_std_logic_vector(2067,16);
	wave(413) <= conv_std_logic_vector(2042,16);
	wave(414) <= conv_std_logic_vector(2035,16);
	wave(415) <= conv_std_logic_vector(2060,16);
	wave(416) <= conv_std_logic_vector(2071,16);
	wave(417) <= conv_std_logic_vector(2048,16);
	wave(418) <= conv_std_logic_vector(2033,16);
	wave(419) <= conv_std_logic_vector(2054,16);
	wave(420) <= conv_std_logic_vector(2072,16);
	wave(421) <= conv_std_logic_vector(2055,16);
	wave(422) <= conv_std_logic_vector(2033,16);
	wave(423) <= conv_std_logic_vector(2047,16);
	wave(424) <= conv_std_logic_vector(2071,16);
	wave(425) <= conv_std_logic_vector(2062,16);
	wave(426) <= conv_std_logic_vector(2037,16);
	wave(427) <= conv_std_logic_vector(2040,16);
	wave(428) <= conv_std_logic_vector(2066,16);
	wave(429) <= conv_std_logic_vector(2069,16);
	wave(430) <= conv_std_logic_vector(2042,16);
	wave(431) <= conv_std_logic_vector(2035,16);
	wave(432) <= conv_std_logic_vector(2061,16);
	wave(433) <= conv_std_logic_vector(2071,16);
	wave(434) <= conv_std_logic_vector(2048,16);
	wave(435) <= conv_std_logic_vector(2034,16);
	wave(436) <= conv_std_logic_vector(2053,16);
	wave(437) <= conv_std_logic_vector(2072,16);
	wave(438) <= conv_std_logic_vector(2057,16);
	wave(439) <= conv_std_logic_vector(2034,16);
	wave(440) <= conv_std_logic_vector(2046,16);
	wave(441) <= conv_std_logic_vector(2070,16);
	wave(442) <= conv_std_logic_vector(2063,16);
	wave(443) <= conv_std_logic_vector(2038,16);
	wave(444) <= conv_std_logic_vector(2039,16);
	wave(445) <= conv_std_logic_vector(2065,16);
	wave(446) <= conv_std_logic_vector(2069,16);
	wave(447) <= conv_std_logic_vector(2043,16);
	wave(448) <= conv_std_logic_vector(2035,16);
	wave(449) <= conv_std_logic_vector(2059,16);
	wave(450) <= conv_std_logic_vector(2072,16);
	wave(451) <= conv_std_logic_vector(2050,16);
	wave(452) <= conv_std_logic_vector(2033,16);
	wave(453) <= conv_std_logic_vector(2052,16);
	wave(454) <= conv_std_logic_vector(2071,16);
	wave(455) <= conv_std_logic_vector(2056,16);
	wave(456) <= conv_std_logic_vector(2034,16);
	wave(457) <= conv_std_logic_vector(2046,16);
	wave(458) <= conv_std_logic_vector(2070,16);
	wave(459) <= conv_std_logic_vector(2063,16);
	wave(460) <= conv_std_logic_vector(2035,16);
	wave(461) <= conv_std_logic_vector(2039,16);
	wave(462) <= conv_std_logic_vector(2068,16);
	wave(463) <= conv_std_logic_vector(2068,16);
	wave(464) <= conv_std_logic_vector(2039,16);
	wave(465) <= conv_std_logic_vector(2036,16);
	wave(466) <= conv_std_logic_vector(2061,16);
	wave(467) <= conv_std_logic_vector(2070,16);
	wave(468) <= conv_std_logic_vector(2045,16);
	wave(469) <= conv_std_logic_vector(2033,16);
	wave(470) <= conv_std_logic_vector(2054,16);
	wave(471) <= conv_std_logic_vector(2070,16);
	wave(472) <= conv_std_logic_vector(2053,16);
	wave(473) <= conv_std_logic_vector(2032,16);
	wave(474) <= conv_std_logic_vector(2047,16);
	wave(475) <= conv_std_logic_vector(2069,16);
	wave(476) <= conv_std_logic_vector(2060,16);
	wave(477) <= conv_std_logic_vector(2032,16);
	wave(478) <= conv_std_logic_vector(2042,16);
	wave(479) <= conv_std_logic_vector(2066,16);
	wave(480) <= conv_std_logic_vector(2066,16);
	wave(481) <= conv_std_logic_vector(2040,16);
	wave(482) <= conv_std_logic_vector(2034,16);
	wave(483) <= conv_std_logic_vector(2058,16);
	wave(484) <= conv_std_logic_vector(2068,16);
	wave(485) <= conv_std_logic_vector(2044,16);
	wave(486) <= conv_std_logic_vector(2032,16);
	wave(487) <= conv_std_logic_vector(2055,16);
	wave(488) <= conv_std_logic_vector(2069,16);
	wave(489) <= conv_std_logic_vector(2050,16);
	wave(490) <= conv_std_logic_vector(2032,16);
	wave(491) <= conv_std_logic_vector(2047,16);
	wave(492) <= conv_std_logic_vector(2068,16);
	wave(493) <= conv_std_logic_vector(2058,16);
	wave(494) <= conv_std_logic_vector(2034,16);
	wave(495) <= conv_std_logic_vector(2039,16);
	wave(496) <= conv_std_logic_vector(2065,16);
	wave(497) <= conv_std_logic_vector(2066,16);
	wave(498) <= conv_std_logic_vector(2038,16);
	wave(499) <= conv_std_logic_vector(2033,16);
	wave(500) <= conv_std_logic_vector(2061,16);
	wave(501) <= conv_std_logic_vector(2061,16);
	wave(502) <= conv_std_logic_vector(2067,16);
	wave(503) <= conv_std_logic_vector(2044,16);
	wave(504) <= conv_std_logic_vector(2031,16);
	wave(505) <= conv_std_logic_vector(2052,16);
	wave(506) <= conv_std_logic_vector(2069,16);
	wave(507) <= conv_std_logic_vector(2052,16);
	wave(508) <= conv_std_logic_vector(2031,16);
	wave(509) <= conv_std_logic_vector(2045,16);
	wave(510) <= conv_std_logic_vector(2068,16);
	wave(511) <= conv_std_logic_vector(2058,16);
	wave(512) <= conv_std_logic_vector(2033,16);
	wave(513) <= conv_std_logic_vector(2039,16);
	wave(514) <= conv_std_logic_vector(2065,16);
	wave(515) <= conv_std_logic_vector(2063,16);
	wave(516) <= conv_std_logic_vector(2038,16);
	wave(517) <= conv_std_logic_vector(2034,16);
	wave(518) <= conv_std_logic_vector(2059,16);
	wave(519) <= conv_std_logic_vector(2068,16);
	wave(520) <= conv_std_logic_vector(2043,16);
	wave(521) <= conv_std_logic_vector(2030,16);
	wave(522) <= conv_std_logic_vector(2054,16);
	wave(523) <= conv_std_logic_vector(2069,16);
	wave(524) <= conv_std_logic_vector(2049,16);
	wave(525) <= conv_std_logic_vector(2030,16);
	wave(526) <= conv_std_logic_vector(2048,16);
	wave(527) <= conv_std_logic_vector(2069,16);
	wave(528) <= conv_std_logic_vector(2056,16);
	wave(529) <= conv_std_logic_vector(2033,16);
	wave(530) <= conv_std_logic_vector(2041,16);
	wave(531) <= conv_std_logic_vector(2065,16);
	wave(532) <= conv_std_logic_vector(2063,16);
	wave(533) <= conv_std_logic_vector(2037,16);
	wave(534) <= conv_std_logic_vector(2034,16);
	wave(535) <= conv_std_logic_vector(2061,16);
	wave(536) <= conv_std_logic_vector(2068,16);
	wave(537) <= conv_std_logic_vector(2044,16);
	wave(538) <= conv_std_logic_vector(2031,16);
	wave(539) <= conv_std_logic_vector(2055,16);
	wave(540) <= conv_std_logic_vector(2070,16);
	wave(541) <= conv_std_logic_vector(2050,16);
	wave(542) <= conv_std_logic_vector(2031,16);
	wave(543) <= conv_std_logic_vector(2048,16);
	wave(544) <= conv_std_logic_vector(2070,16);
	wave(545) <= conv_std_logic_vector(2057,16);
	wave(546) <= conv_std_logic_vector(2033,16);
	wave(547) <= conv_std_logic_vector(2041,16);
	wave(548) <= conv_std_logic_vector(2065,16);
	wave(549) <= conv_std_logic_vector(2063,16);
	wave(550) <= conv_std_logic_vector(2038,16);
	wave(551) <= conv_std_logic_vector(2037,16);
	wave(552) <= conv_std_logic_vector(2059,16);
	wave(553) <= conv_std_logic_vector(2065,16);
	wave(554) <= conv_std_logic_vector(2046,16);
	wave(555) <= conv_std_logic_vector(2033,16);
	wave(556) <= conv_std_logic_vector(2051,16);
	wave(557) <= conv_std_logic_vector(2069,16);
	wave(558) <= conv_std_logic_vector(2053,16);
	wave(559) <= conv_std_logic_vector(2032,16);
	wave(560) <= conv_std_logic_vector(2044,16);
	wave(561) <= conv_std_logic_vector(2068,16);
	wave(562) <= conv_std_logic_vector(2061,16);
	wave(563) <= conv_std_logic_vector(2034,16);
	wave(564) <= conv_std_logic_vector(2037,16);
	wave(565) <= conv_std_logic_vector(2064,16);
	wave(566) <= conv_std_logic_vector(2065,16);
	wave(567) <= conv_std_logic_vector(2040,16);
	wave(568) <= conv_std_logic_vector(2034,16);
	wave(569) <= conv_std_logic_vector(2054,16);
	wave(570) <= conv_std_logic_vector(2067,16);
	wave(571) <= conv_std_logic_vector(2046,16);
	wave(572) <= conv_std_logic_vector(2030,16);
	wave(573) <= conv_std_logic_vector(2052,16);
	wave(574) <= conv_std_logic_vector(2069,16);
	wave(575) <= conv_std_logic_vector(2049,16);
	wave(576) <= conv_std_logic_vector(2030,16);
	wave(577) <= conv_std_logic_vector(2046,16);
	wave(578) <= conv_std_logic_vector(2066,16);
	wave(579) <= conv_std_logic_vector(2057,16);
	wave(580) <= conv_std_logic_vector(2033,16);
	wave(581) <= conv_std_logic_vector(2038,16);
	wave(582) <= conv_std_logic_vector(2063,16);
	wave(583) <= conv_std_logic_vector(2064,16);
	wave(584) <= conv_std_logic_vector(2037,16);
	wave(585) <= conv_std_logic_vector(2032,16);
	wave(586) <= conv_std_logic_vector(2058,16);
	wave(587) <= conv_std_logic_vector(2067,16);
	wave(588) <= conv_std_logic_vector(2044,16);
	wave(589) <= conv_std_logic_vector(2029,16);
	wave(590) <= conv_std_logic_vector(2050,16);
	wave(591) <= conv_std_logic_vector(2068,16);
	wave(592) <= conv_std_logic_vector(2050,16);
	wave(593) <= conv_std_logic_vector(2029,16);
	wave(594) <= conv_std_logic_vector(2044,16);
	wave(595) <= conv_std_logic_vector(2066,16);
	wave(596) <= conv_std_logic_vector(2057,16);
	wave(597) <= conv_std_logic_vector(2031,16);
	wave(598) <= conv_std_logic_vector(2037,16);
	wave(599) <= conv_std_logic_vector(2064,16);
	wave(600) <= conv_std_logic_vector(2062,16);
	wave(601) <= conv_std_logic_vector(2036,16);
	wave(602) <= conv_std_logic_vector(2033,16);
	wave(603) <= conv_std_logic_vector(2059,16);
	wave(604) <= conv_std_logic_vector(2066,16);
	wave(605) <= conv_std_logic_vector(2042,16);
	wave(606) <= conv_std_logic_vector(2029,16);
	wave(607) <= conv_std_logic_vector(2053,16);
	wave(608) <= conv_std_logic_vector(2067,16);
	wave(609) <= conv_std_logic_vector(2047,16);
	wave(610) <= conv_std_logic_vector(2030,16);
	wave(611) <= conv_std_logic_vector(2046,16);
	wave(612) <= conv_std_logic_vector(2068,16);
	wave(613) <= conv_std_logic_vector(2053,16);
	wave(614) <= conv_std_logic_vector(2030,16);
	wave(615) <= conv_std_logic_vector(2040,16);
	wave(616) <= conv_std_logic_vector(2065,16);
	wave(617) <= conv_std_logic_vector(2059,16);
	wave(618) <= conv_std_logic_vector(2033,16);
	wave(619) <= conv_std_logic_vector(2035,16);
	wave(620) <= conv_std_logic_vector(2061,16);
	wave(621) <= conv_std_logic_vector(2066,16);
	wave(622) <= conv_std_logic_vector(2038,16);
	wave(623) <= conv_std_logic_vector(2031,16);
	wave(624) <= conv_std_logic_vector(2056,16);
	wave(625) <= conv_std_logic_vector(2067,16);
	wave(626) <= conv_std_logic_vector(2043,16);
	wave(627) <= conv_std_logic_vector(2028,16);
	wave(628) <= conv_std_logic_vector(2051,16);
	wave(629) <= conv_std_logic_vector(2068,16);
	wave(630) <= conv_std_logic_vector(2049,16);
	wave(631) <= conv_std_logic_vector(2029,16);
	wave(632) <= conv_std_logic_vector(2044,16);
	wave(633) <= conv_std_logic_vector(2065,16);
	wave(634) <= conv_std_logic_vector(2057,16);
	wave(635) <= conv_std_logic_vector(2032,16);
	wave(636) <= conv_std_logic_vector(2036,16);
	wave(637) <= conv_std_logic_vector(2062,16);
	wave(638) <= conv_std_logic_vector(2063,16);
	wave(639) <= conv_std_logic_vector(2036,16);
	wave(640) <= conv_std_logic_vector(2030,16);
	wave(641) <= conv_std_logic_vector(2058,16);
	wave(642) <= conv_std_logic_vector(2069,16);
	wave(643) <= conv_std_logic_vector(2041,16);
	wave(644) <= conv_std_logic_vector(2027,16);
	wave(645) <= conv_std_logic_vector(2052,16);
	wave(646) <= conv_std_logic_vector(2069,16);
	wave(647) <= conv_std_logic_vector(2049,16);
	wave(648) <= conv_std_logic_vector(2028,16);
	wave(649) <= conv_std_logic_vector(2045,16);
	wave(650) <= conv_std_logic_vector(2065,16);
	wave(651) <= conv_std_logic_vector(2056,16);
	wave(652) <= conv_std_logic_vector(2033,16);
	wave(653) <= conv_std_logic_vector(2035,16);
	wave(654) <= conv_std_logic_vector(2059,16);
	wave(655) <= conv_std_logic_vector(2064,16);
	wave(656) <= conv_std_logic_vector(2038,16);
	wave(657) <= conv_std_logic_vector(2030,16);
	wave(658) <= conv_std_logic_vector(2058,16);
	wave(659) <= conv_std_logic_vector(2067,16);
	wave(660) <= conv_std_logic_vector(2044,16);
	wave(661) <= conv_std_logic_vector(2028,16);
	wave(662) <= conv_std_logic_vector(2047,16);
	wave(663) <= conv_std_logic_vector(2066,16);
	wave(664) <= conv_std_logic_vector(2051,16);
	wave(665) <= conv_std_logic_vector(2027,16);
	wave(666) <= conv_std_logic_vector(2042,16);
	wave(667) <= conv_std_logic_vector(2065,16);
	wave(668) <= conv_std_logic_vector(2057,16);
	wave(669) <= conv_std_logic_vector(2030,16);
	wave(670) <= conv_std_logic_vector(2035,16);
	wave(671) <= conv_std_logic_vector(2062,16);
	wave(672) <= conv_std_logic_vector(2063,16);
	wave(673) <= conv_std_logic_vector(2035,16);
	wave(674) <= conv_std_logic_vector(2030,16);
	wave(675) <= conv_std_logic_vector(2056,16);
	wave(676) <= conv_std_logic_vector(2065,16);
	wave(677) <= conv_std_logic_vector(2040,16);
	wave(678) <= conv_std_logic_vector(2028,16);
	wave(679) <= conv_std_logic_vector(2051,16);
	wave(680) <= conv_std_logic_vector(2066,16);
	wave(681) <= conv_std_logic_vector(2046,16);
	wave(682) <= conv_std_logic_vector(2027,16);
	wave(683) <= conv_std_logic_vector(2043,16);
	wave(684) <= conv_std_logic_vector(2066,16);
	wave(685) <= conv_std_logic_vector(2053,16);
	wave(686) <= conv_std_logic_vector(2028,16);
	wave(687) <= conv_std_logic_vector(2037,16);
	wave(688) <= conv_std_logic_vector(2062,16);
	wave(689) <= conv_std_logic_vector(2060,16);
	wave(690) <= conv_std_logic_vector(2033,16);
	wave(691) <= conv_std_logic_vector(2030,16);
	wave(692) <= conv_std_logic_vector(2056,16);
	wave(693) <= conv_std_logic_vector(2064,16);
	wave(694) <= conv_std_logic_vector(2039,16);
	wave(695) <= conv_std_logic_vector(2028,16);
	wave(696) <= conv_std_logic_vector(2051,16);
	wave(697) <= conv_std_logic_vector(2066,16);
	wave(698) <= conv_std_logic_vector(2046,16);
	wave(699) <= conv_std_logic_vector(2026,16);
	wave(700) <= conv_std_logic_vector(2045,16);
	wave(701) <= conv_std_logic_vector(2066,16);
	wave(702) <= conv_std_logic_vector(2052,16);
	wave(703) <= conv_std_logic_vector(2028,16);
	wave(704) <= conv_std_logic_vector(2040,16);
	wave(705) <= conv_std_logic_vector(2065,16);
	wave(706) <= conv_std_logic_vector(2058,16);
	wave(707) <= conv_std_logic_vector(2032,16);
	wave(708) <= conv_std_logic_vector(2034,16);
	wave(709) <= conv_std_logic_vector(2060,16);
	wave(710) <= conv_std_logic_vector(2064,16);
	wave(711) <= conv_std_logic_vector(2038,16);
	wave(712) <= conv_std_logic_vector(2030,16);
	wave(713) <= conv_std_logic_vector(2055,16);
	wave(714) <= conv_std_logic_vector(2067,16);
	wave(715) <= conv_std_logic_vector(2044,16);
	wave(716) <= conv_std_logic_vector(2028,16);
	wave(717) <= conv_std_logic_vector(2049,16);
	wave(718) <= conv_std_logic_vector(2067,16);
	wave(719) <= conv_std_logic_vector(2051,16);
	wave(720) <= conv_std_logic_vector(2028,16);
	wave(721) <= conv_std_logic_vector(2042,16);
	wave(722) <= conv_std_logic_vector(2066,16);
	wave(723) <= conv_std_logic_vector(2057,16);
	wave(724) <= conv_std_logic_vector(2032,16);
	wave(725) <= conv_std_logic_vector(2036,16);
	wave(726) <= conv_std_logic_vector(2062,16);
	wave(727) <= conv_std_logic_vector(2063,16);
	wave(728) <= conv_std_logic_vector(2037,16);
	wave(729) <= conv_std_logic_vector(2032,16);
	wave(730) <= conv_std_logic_vector(2059,16);
	wave(731) <= conv_std_logic_vector(2064,16);
	wave(732) <= conv_std_logic_vector(2040,16);
	wave(733) <= conv_std_logic_vector(2030,16);
	wave(734) <= conv_std_logic_vector(2053,16);
	wave(735) <= conv_std_logic_vector(2067,16);
	wave(736) <= conv_std_logic_vector(2047,16);
	wave(737) <= conv_std_logic_vector(2028,16);
	wave(738) <= conv_std_logic_vector(2048,16);
	wave(739) <= conv_std_logic_vector(2067,16);
	wave(740) <= conv_std_logic_vector(2052,16);
	wave(741) <= conv_std_logic_vector(2029,16);
	wave(742) <= conv_std_logic_vector(2042,16);
	wave(743) <= conv_std_logic_vector(2066,16);
	wave(744) <= conv_std_logic_vector(2058,16);
	wave(745) <= conv_std_logic_vector(2032,16);
	wave(746) <= conv_std_logic_vector(2036,16);
	wave(747) <= conv_std_logic_vector(2060,16);
	wave(748) <= conv_std_logic_vector(2062,16);
	wave(749) <= conv_std_logic_vector(2035,16);
	wave(750) <= conv_std_logic_vector(2032,16);
	wave(751) <= conv_std_logic_vector(2061,16);
	wave(752) <= conv_std_logic_vector(2067,16);
	wave(753) <= conv_std_logic_vector(2040,16);
	wave(754) <= conv_std_logic_vector(2028,16);
	wave(755) <= conv_std_logic_vector(2055,16);
	wave(756) <= conv_std_logic_vector(2068,16);
	wave(757) <= conv_std_logic_vector(2045,16);
	wave(758) <= conv_std_logic_vector(2028,16);
	wave(759) <= conv_std_logic_vector(2048,16);
	wave(760) <= conv_std_logic_vector(2067,16);
	wave(761) <= conv_std_logic_vector(2051,16);
	wave(762) <= conv_std_logic_vector(2028,16);
	wave(763) <= conv_std_logic_vector(2042,16);
	wave(764) <= conv_std_logic_vector(2066,16);
	wave(765) <= conv_std_logic_vector(2056,16);
	wave(766) <= conv_std_logic_vector(2028,16);
	wave(767) <= conv_std_logic_vector(2037,16);

end Behavioral;